// nios_sys.v

// Generated using ACDS version 13.0sp1 232 at 2025.04.25.22:56:28

`timescale 1 ps / 1 ps
module nios_sys (
		input  wire       clk_clk,                             //                          clk.clk
		input  wire       reset_reset_n,                       //                        reset.reset_n
		output wire [7:0] lcd_data_external_connection_export, // lcd_data_external_connection.export
		output wire       lcd_rw_external_connection_export,   //   lcd_rw_external_connection.export
		output wire       lcd_rs_external_connection_export,   //   lcd_rs_external_connection.export
		output wire       lcd_en_external_connection_export,   //   lcd_en_external_connection.export
		output wire       lcd_on_external_connection_export,   //   lcd_on_external_connection.export
		output wire [7:0] led8_external_connection_export,     //     led8_external_connection.export
		output wire [7:0] led7_external_connection_export,     //     led7_external_connection.export
		output wire [7:0] led6_external_connection_export,     //     led6_external_connection.export
		output wire [7:0] led5_external_connection_export,     //     led5_external_connection.export
		output wire [7:0] led4_external_connection_export,     //     led4_external_connection.export
		output wire [7:0] led3_external_connection_export,     //     led3_external_connection.export
		output wire [7:0] led2_external_connection_export,     //     led2_external_connection.export
		output wire [7:0] led1_external_connection_export,     //     led1_external_connection.export
		input  wire       uart_0_external_connection_rxd,      //   uart_0_external_connection.rxd
		output wire       uart_0_external_connection_txd,      //                             .txd
		input  wire [1:0] switch0_external_connection_export,  //  switch0_external_connection.export
		input  wire       key3_external_connection_export,     //     key3_external_connection.export
		input  wire       key2_external_connection_export,     //     key2_external_connection.export
		input  wire       key1_external_connection_export,     //     key1_external_connection.export
		output wire [7:0] ledr_external_connection_export      //     ledr_external_connection.export
	);

	wire         nios2_qsys_0_instruction_master_waitrequest;                                                         // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [20:0] nios2_qsys_0_instruction_master_address;                                                             // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire         nios2_qsys_0_instruction_master_read;                                                                // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                                            // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                                                // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                                                  // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire  [20:0] nios2_qsys_0_data_master_address;                                                                    // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire         nios2_qsys_0_data_master_write;                                                                      // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire         nios2_qsys_0_data_master_read;                                                                       // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                                                   // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                                                // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                                                 // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                           // nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                  // nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                        // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire  [16:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                          // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                       // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                            // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                            // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                         // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                       // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [31:0] led8_s1_translator_avalon_anti_slave_0_writedata;                                                    // led8_s1_translator:av_writedata -> led8:writedata
	wire   [1:0] led8_s1_translator_avalon_anti_slave_0_address;                                                      // led8_s1_translator:av_address -> led8:address
	wire         led8_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led8_s1_translator:av_chipselect -> led8:chipselect
	wire         led8_s1_translator_avalon_anti_slave_0_write;                                                        // led8_s1_translator:av_write -> led8:write_n
	wire  [31:0] led8_s1_translator_avalon_anti_slave_0_readdata;                                                     // led8:readdata -> led8_s1_translator:av_readdata
	wire  [31:0] led7_s1_translator_avalon_anti_slave_0_writedata;                                                    // led7_s1_translator:av_writedata -> led7:writedata
	wire   [1:0] led7_s1_translator_avalon_anti_slave_0_address;                                                      // led7_s1_translator:av_address -> led7:address
	wire         led7_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led7_s1_translator:av_chipselect -> led7:chipselect
	wire         led7_s1_translator_avalon_anti_slave_0_write;                                                        // led7_s1_translator:av_write -> led7:write_n
	wire  [31:0] led7_s1_translator_avalon_anti_slave_0_readdata;                                                     // led7:readdata -> led7_s1_translator:av_readdata
	wire  [31:0] led6_s1_translator_avalon_anti_slave_0_writedata;                                                    // led6_s1_translator:av_writedata -> led6:writedata
	wire   [1:0] led6_s1_translator_avalon_anti_slave_0_address;                                                      // led6_s1_translator:av_address -> led6:address
	wire         led6_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led6_s1_translator:av_chipselect -> led6:chipselect
	wire         led6_s1_translator_avalon_anti_slave_0_write;                                                        // led6_s1_translator:av_write -> led6:write_n
	wire  [31:0] led6_s1_translator_avalon_anti_slave_0_readdata;                                                     // led6:readdata -> led6_s1_translator:av_readdata
	wire  [31:0] led5_s1_translator_avalon_anti_slave_0_writedata;                                                    // led5_s1_translator:av_writedata -> led5:writedata
	wire   [1:0] led5_s1_translator_avalon_anti_slave_0_address;                                                      // led5_s1_translator:av_address -> led5:address
	wire         led5_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led5_s1_translator:av_chipselect -> led5:chipselect
	wire         led5_s1_translator_avalon_anti_slave_0_write;                                                        // led5_s1_translator:av_write -> led5:write_n
	wire  [31:0] led5_s1_translator_avalon_anti_slave_0_readdata;                                                     // led5:readdata -> led5_s1_translator:av_readdata
	wire  [31:0] led4_s1_translator_avalon_anti_slave_0_writedata;                                                    // led4_s1_translator:av_writedata -> led4:writedata
	wire   [1:0] led4_s1_translator_avalon_anti_slave_0_address;                                                      // led4_s1_translator:av_address -> led4:address
	wire         led4_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led4_s1_translator:av_chipselect -> led4:chipselect
	wire         led4_s1_translator_avalon_anti_slave_0_write;                                                        // led4_s1_translator:av_write -> led4:write_n
	wire  [31:0] led4_s1_translator_avalon_anti_slave_0_readdata;                                                     // led4:readdata -> led4_s1_translator:av_readdata
	wire  [31:0] led3_s1_translator_avalon_anti_slave_0_writedata;                                                    // led3_s1_translator:av_writedata -> led3:writedata
	wire   [1:0] led3_s1_translator_avalon_anti_slave_0_address;                                                      // led3_s1_translator:av_address -> led3:address
	wire         led3_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led3_s1_translator:av_chipselect -> led3:chipselect
	wire         led3_s1_translator_avalon_anti_slave_0_write;                                                        // led3_s1_translator:av_write -> led3:write_n
	wire  [31:0] led3_s1_translator_avalon_anti_slave_0_readdata;                                                     // led3:readdata -> led3_s1_translator:av_readdata
	wire  [31:0] led2_s1_translator_avalon_anti_slave_0_writedata;                                                    // led2_s1_translator:av_writedata -> led2:writedata
	wire   [1:0] led2_s1_translator_avalon_anti_slave_0_address;                                                      // led2_s1_translator:av_address -> led2:address
	wire         led2_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led2_s1_translator:av_chipselect -> led2:chipselect
	wire         led2_s1_translator_avalon_anti_slave_0_write;                                                        // led2_s1_translator:av_write -> led2:write_n
	wire  [31:0] led2_s1_translator_avalon_anti_slave_0_readdata;                                                     // led2:readdata -> led2_s1_translator:av_readdata
	wire  [31:0] led1_s1_translator_avalon_anti_slave_0_writedata;                                                    // led1_s1_translator:av_writedata -> led1:writedata
	wire   [1:0] led1_s1_translator_avalon_anti_slave_0_address;                                                      // led1_s1_translator:av_address -> led1:address
	wire         led1_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led1_s1_translator:av_chipselect -> led1:chipselect
	wire         led1_s1_translator_avalon_anti_slave_0_write;                                                        // led1_s1_translator:av_write -> led1:write_n
	wire  [31:0] led1_s1_translator_avalon_anti_slave_0_readdata;                                                     // led1:readdata -> led1_s1_translator:av_readdata
	wire  [15:0] uart_0_s1_translator_avalon_anti_slave_0_writedata;                                                  // uart_0_s1_translator:av_writedata -> uart_0:writedata
	wire   [2:0] uart_0_s1_translator_avalon_anti_slave_0_address;                                                    // uart_0_s1_translator:av_address -> uart_0:address
	wire         uart_0_s1_translator_avalon_anti_slave_0_chipselect;                                                 // uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	wire         uart_0_s1_translator_avalon_anti_slave_0_write;                                                      // uart_0_s1_translator:av_write -> uart_0:write_n
	wire         uart_0_s1_translator_avalon_anti_slave_0_read;                                                       // uart_0_s1_translator:av_read -> uart_0:read_n
	wire  [15:0] uart_0_s1_translator_avalon_anti_slave_0_readdata;                                                   // uart_0:readdata -> uart_0_s1_translator:av_readdata
	wire         uart_0_s1_translator_avalon_anti_slave_0_begintransfer;                                              // uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	wire  [31:0] switch0_s1_translator_avalon_anti_slave_0_writedata;                                                 // switch0_s1_translator:av_writedata -> switch0:writedata
	wire   [1:0] switch0_s1_translator_avalon_anti_slave_0_address;                                                   // switch0_s1_translator:av_address -> switch0:address
	wire         switch0_s1_translator_avalon_anti_slave_0_chipselect;                                                // switch0_s1_translator:av_chipselect -> switch0:chipselect
	wire         switch0_s1_translator_avalon_anti_slave_0_write;                                                     // switch0_s1_translator:av_write -> switch0:write_n
	wire  [31:0] switch0_s1_translator_avalon_anti_slave_0_readdata;                                                  // switch0:readdata -> switch0_s1_translator:av_readdata
	wire   [1:0] key3_s1_translator_avalon_anti_slave_0_address;                                                      // key3_s1_translator:av_address -> key3:address
	wire  [31:0] key3_s1_translator_avalon_anti_slave_0_readdata;                                                     // key3:readdata -> key3_s1_translator:av_readdata
	wire   [1:0] key2_s1_translator_avalon_anti_slave_0_address;                                                      // key2_s1_translator:av_address -> key2:address
	wire  [31:0] key2_s1_translator_avalon_anti_slave_0_readdata;                                                     // key2:readdata -> key2_s1_translator:av_readdata
	wire   [1:0] key1_s1_translator_avalon_anti_slave_0_address;                                                      // key1_s1_translator:av_address -> key1:address
	wire  [31:0] key1_s1_translator_avalon_anti_slave_0_readdata;                                                     // key1:readdata -> key1_s1_translator:av_readdata
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                   // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                     // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire  [31:0] ledr_s1_translator_avalon_anti_slave_0_writedata;                                                    // ledr_s1_translator:av_writedata -> ledr:writedata
	wire   [1:0] ledr_s1_translator_avalon_anti_slave_0_address;                                                      // ledr_s1_translator:av_address -> ledr:address
	wire         ledr_s1_translator_avalon_anti_slave_0_chipselect;                                                   // ledr_s1_translator:av_chipselect -> ledr:chipselect
	wire         ledr_s1_translator_avalon_anti_slave_0_write;                                                        // ledr_s1_translator:av_write -> ledr:write_n
	wire  [31:0] ledr_s1_translator_avalon_anti_slave_0_readdata;                                                     // ledr:readdata -> ledr_s1_translator:av_readdata
	wire  [31:0] lcd_data_s1_translator_avalon_anti_slave_0_writedata;                                                // LCD_DATA_s1_translator:av_writedata -> LCD_DATA:writedata
	wire   [1:0] lcd_data_s1_translator_avalon_anti_slave_0_address;                                                  // LCD_DATA_s1_translator:av_address -> LCD_DATA:address
	wire         lcd_data_s1_translator_avalon_anti_slave_0_chipselect;                                               // LCD_DATA_s1_translator:av_chipselect -> LCD_DATA:chipselect
	wire         lcd_data_s1_translator_avalon_anti_slave_0_write;                                                    // LCD_DATA_s1_translator:av_write -> LCD_DATA:write_n
	wire  [31:0] lcd_data_s1_translator_avalon_anti_slave_0_readdata;                                                 // LCD_DATA:readdata -> LCD_DATA_s1_translator:av_readdata
	wire  [31:0] lcd_rw_s1_translator_avalon_anti_slave_0_writedata;                                                  // LCD_RW_s1_translator:av_writedata -> LCD_RW:writedata
	wire   [1:0] lcd_rw_s1_translator_avalon_anti_slave_0_address;                                                    // LCD_RW_s1_translator:av_address -> LCD_RW:address
	wire         lcd_rw_s1_translator_avalon_anti_slave_0_chipselect;                                                 // LCD_RW_s1_translator:av_chipselect -> LCD_RW:chipselect
	wire         lcd_rw_s1_translator_avalon_anti_slave_0_write;                                                      // LCD_RW_s1_translator:av_write -> LCD_RW:write_n
	wire  [31:0] lcd_rw_s1_translator_avalon_anti_slave_0_readdata;                                                   // LCD_RW:readdata -> LCD_RW_s1_translator:av_readdata
	wire  [31:0] lcd_rs_s1_translator_avalon_anti_slave_0_writedata;                                                  // LCD_RS_s1_translator:av_writedata -> LCD_RS:writedata
	wire   [1:0] lcd_rs_s1_translator_avalon_anti_slave_0_address;                                                    // LCD_RS_s1_translator:av_address -> LCD_RS:address
	wire         lcd_rs_s1_translator_avalon_anti_slave_0_chipselect;                                                 // LCD_RS_s1_translator:av_chipselect -> LCD_RS:chipselect
	wire         lcd_rs_s1_translator_avalon_anti_slave_0_write;                                                      // LCD_RS_s1_translator:av_write -> LCD_RS:write_n
	wire  [31:0] lcd_rs_s1_translator_avalon_anti_slave_0_readdata;                                                   // LCD_RS:readdata -> LCD_RS_s1_translator:av_readdata
	wire  [31:0] lcd_en_s1_translator_avalon_anti_slave_0_writedata;                                                  // LCD_EN_s1_translator:av_writedata -> LCD_EN:writedata
	wire   [1:0] lcd_en_s1_translator_avalon_anti_slave_0_address;                                                    // LCD_EN_s1_translator:av_address -> LCD_EN:address
	wire         lcd_en_s1_translator_avalon_anti_slave_0_chipselect;                                                 // LCD_EN_s1_translator:av_chipselect -> LCD_EN:chipselect
	wire         lcd_en_s1_translator_avalon_anti_slave_0_write;                                                      // LCD_EN_s1_translator:av_write -> LCD_EN:write_n
	wire  [31:0] lcd_en_s1_translator_avalon_anti_slave_0_readdata;                                                   // LCD_EN:readdata -> LCD_EN_s1_translator:av_readdata
	wire  [31:0] lcd_on_s1_translator_avalon_anti_slave_0_writedata;                                                  // LCD_ON_s1_translator:av_writedata -> LCD_ON:writedata
	wire   [1:0] lcd_on_s1_translator_avalon_anti_slave_0_address;                                                    // LCD_ON_s1_translator:av_address -> LCD_ON:address
	wire         lcd_on_s1_translator_avalon_anti_slave_0_chipselect;                                                 // LCD_ON_s1_translator:av_chipselect -> LCD_ON:chipselect
	wire         lcd_on_s1_translator_avalon_anti_slave_0_write;                                                      // LCD_ON_s1_translator:av_write -> LCD_ON:write_n
	wire  [31:0] lcd_on_s1_translator_avalon_anti_slave_0_readdata;                                                   // LCD_ON:readdata -> LCD_ON_s1_translator:av_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire  [20:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire  [20:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [20:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led8_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led8_s1_translator:uav_waitrequest -> led8_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led8_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led8_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led8_s1_translator:uav_burstcount
	wire  [31:0] led8_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led8_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led8_s1_translator:uav_writedata
	wire  [20:0] led8_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led8_s1_translator_avalon_universal_slave_0_agent:m0_address -> led8_s1_translator:uav_address
	wire         led8_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led8_s1_translator_avalon_universal_slave_0_agent:m0_write -> led8_s1_translator:uav_write
	wire         led8_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led8_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led8_s1_translator:uav_lock
	wire         led8_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led8_s1_translator_avalon_universal_slave_0_agent:m0_read -> led8_s1_translator:uav_read
	wire  [31:0] led8_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led8_s1_translator:uav_readdata -> led8_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led8_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led8_s1_translator:uav_readdatavalid -> led8_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led8_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led8_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led8_s1_translator:uav_debugaccess
	wire   [3:0] led8_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led8_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led8_s1_translator:uav_byteenable
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led8_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led8_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led8_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led8_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led8_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led8_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led8_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led8_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led8_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led8_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led8_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led7_s1_translator:uav_waitrequest -> led7_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led7_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led7_s1_translator:uav_burstcount
	wire  [31:0] led7_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led7_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led7_s1_translator:uav_writedata
	wire  [20:0] led7_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led7_s1_translator_avalon_universal_slave_0_agent:m0_address -> led7_s1_translator:uav_address
	wire         led7_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led7_s1_translator_avalon_universal_slave_0_agent:m0_write -> led7_s1_translator:uav_write
	wire         led7_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led7_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led7_s1_translator:uav_lock
	wire         led7_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led7_s1_translator_avalon_universal_slave_0_agent:m0_read -> led7_s1_translator:uav_read
	wire  [31:0] led7_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led7_s1_translator:uav_readdata -> led7_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led7_s1_translator:uav_readdatavalid -> led7_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led7_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led7_s1_translator:uav_debugaccess
	wire   [3:0] led7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led7_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led7_s1_translator:uav_byteenable
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led7_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led7_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led7_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led7_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led7_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led7_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led7_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led7_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led7_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led7_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led7_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led6_s1_translator:uav_waitrequest -> led6_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led6_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led6_s1_translator:uav_burstcount
	wire  [31:0] led6_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led6_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led6_s1_translator:uav_writedata
	wire  [20:0] led6_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led6_s1_translator_avalon_universal_slave_0_agent:m0_address -> led6_s1_translator:uav_address
	wire         led6_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led6_s1_translator_avalon_universal_slave_0_agent:m0_write -> led6_s1_translator:uav_write
	wire         led6_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led6_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led6_s1_translator:uav_lock
	wire         led6_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led6_s1_translator_avalon_universal_slave_0_agent:m0_read -> led6_s1_translator:uav_read
	wire  [31:0] led6_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led6_s1_translator:uav_readdata -> led6_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led6_s1_translator:uav_readdatavalid -> led6_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led6_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led6_s1_translator:uav_debugaccess
	wire   [3:0] led6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led6_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led6_s1_translator:uav_byteenable
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led6_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led6_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led6_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led6_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led6_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led6_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led6_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led6_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led6_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led6_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led6_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led5_s1_translator:uav_waitrequest -> led5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led5_s1_translator:uav_burstcount
	wire  [31:0] led5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led5_s1_translator:uav_writedata
	wire  [20:0] led5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led5_s1_translator_avalon_universal_slave_0_agent:m0_address -> led5_s1_translator:uav_address
	wire         led5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led5_s1_translator_avalon_universal_slave_0_agent:m0_write -> led5_s1_translator:uav_write
	wire         led5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led5_s1_translator:uav_lock
	wire         led5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led5_s1_translator_avalon_universal_slave_0_agent:m0_read -> led5_s1_translator:uav_read
	wire  [31:0] led5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led5_s1_translator:uav_readdata -> led5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led5_s1_translator:uav_readdatavalid -> led5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led5_s1_translator:uav_debugaccess
	wire   [3:0] led5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led5_s1_translator:uav_byteenable
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led4_s1_translator:uav_waitrequest -> led4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led4_s1_translator:uav_burstcount
	wire  [31:0] led4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led4_s1_translator:uav_writedata
	wire  [20:0] led4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led4_s1_translator_avalon_universal_slave_0_agent:m0_address -> led4_s1_translator:uav_address
	wire         led4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led4_s1_translator_avalon_universal_slave_0_agent:m0_write -> led4_s1_translator:uav_write
	wire         led4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led4_s1_translator:uav_lock
	wire         led4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led4_s1_translator_avalon_universal_slave_0_agent:m0_read -> led4_s1_translator:uav_read
	wire  [31:0] led4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led4_s1_translator:uav_readdata -> led4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led4_s1_translator:uav_readdatavalid -> led4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led4_s1_translator:uav_debugaccess
	wire   [3:0] led4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led4_s1_translator:uav_byteenable
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led3_s1_translator:uav_waitrequest -> led3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led3_s1_translator:uav_burstcount
	wire  [31:0] led3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led3_s1_translator:uav_writedata
	wire  [20:0] led3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led3_s1_translator_avalon_universal_slave_0_agent:m0_address -> led3_s1_translator:uav_address
	wire         led3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led3_s1_translator_avalon_universal_slave_0_agent:m0_write -> led3_s1_translator:uav_write
	wire         led3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led3_s1_translator:uav_lock
	wire         led3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led3_s1_translator_avalon_universal_slave_0_agent:m0_read -> led3_s1_translator:uav_read
	wire  [31:0] led3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led3_s1_translator:uav_readdata -> led3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led3_s1_translator:uav_readdatavalid -> led3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led3_s1_translator:uav_debugaccess
	wire   [3:0] led3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led3_s1_translator:uav_byteenable
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led2_s1_translator:uav_waitrequest -> led2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led2_s1_translator:uav_burstcount
	wire  [31:0] led2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led2_s1_translator:uav_writedata
	wire  [20:0] led2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led2_s1_translator_avalon_universal_slave_0_agent:m0_address -> led2_s1_translator:uav_address
	wire         led2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led2_s1_translator_avalon_universal_slave_0_agent:m0_write -> led2_s1_translator:uav_write
	wire         led2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led2_s1_translator:uav_lock
	wire         led2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led2_s1_translator_avalon_universal_slave_0_agent:m0_read -> led2_s1_translator:uav_read
	wire  [31:0] led2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led2_s1_translator:uav_readdata -> led2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led2_s1_translator:uav_readdatavalid -> led2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led2_s1_translator:uav_debugaccess
	wire   [3:0] led2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led2_s1_translator:uav_byteenable
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led1_s1_translator:uav_waitrequest -> led1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led1_s1_translator:uav_burstcount
	wire  [31:0] led1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led1_s1_translator:uav_writedata
	wire  [20:0] led1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led1_s1_translator_avalon_universal_slave_0_agent:m0_address -> led1_s1_translator:uav_address
	wire         led1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led1_s1_translator_avalon_universal_slave_0_agent:m0_write -> led1_s1_translator:uav_write
	wire         led1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led1_s1_translator:uav_lock
	wire         led1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led1_s1_translator_avalon_universal_slave_0_agent:m0_read -> led1_s1_translator:uav_read
	wire  [31:0] led1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led1_s1_translator:uav_readdata -> led1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led1_s1_translator:uav_readdatavalid -> led1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led1_s1_translator:uav_debugaccess
	wire   [3:0] led1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led1_s1_translator:uav_byteenable
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] led1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // uart_0_s1_translator:uav_waitrequest -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_0_s1_translator:uav_burstcount
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_0_s1_translator:uav_writedata
	wire  [20:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_0_s1_translator:uav_address
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_0_s1_translator:uav_write
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_0_s1_translator:uav_lock
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_0_s1_translator:uav_read
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // uart_0_s1_translator:uav_readdata -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // uart_0_s1_translator:uav_readdatavalid -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_0_s1_translator:uav_debugaccess
	wire   [3:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_0_s1_translator:uav_byteenable
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // switch0_s1_translator:uav_waitrequest -> switch0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // switch0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch0_s1_translator:uav_burstcount
	wire  [31:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // switch0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch0_s1_translator:uav_writedata
	wire  [20:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // switch0_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch0_s1_translator:uav_address
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // switch0_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch0_s1_translator:uav_write
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // switch0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch0_s1_translator:uav_lock
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // switch0_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch0_s1_translator:uav_read
	wire  [31:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // switch0_s1_translator:uav_readdata -> switch0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // switch0_s1_translator:uav_readdatavalid -> switch0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // switch0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch0_s1_translator:uav_debugaccess
	wire   [3:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // switch0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch0_s1_translator:uav_byteenable
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // key3_s1_translator:uav_waitrequest -> key3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // key3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key3_s1_translator:uav_burstcount
	wire  [31:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // key3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key3_s1_translator:uav_writedata
	wire  [20:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // key3_s1_translator_avalon_universal_slave_0_agent:m0_address -> key3_s1_translator:uav_address
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // key3_s1_translator_avalon_universal_slave_0_agent:m0_write -> key3_s1_translator:uav_write
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // key3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key3_s1_translator:uav_lock
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // key3_s1_translator_avalon_universal_slave_0_agent:m0_read -> key3_s1_translator:uav_read
	wire  [31:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // key3_s1_translator:uav_readdata -> key3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // key3_s1_translator:uav_readdatavalid -> key3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // key3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key3_s1_translator:uav_debugaccess
	wire   [3:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // key3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key3_s1_translator:uav_byteenable
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] key3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // key2_s1_translator:uav_waitrequest -> key2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // key2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key2_s1_translator:uav_burstcount
	wire  [31:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // key2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key2_s1_translator:uav_writedata
	wire  [20:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // key2_s1_translator_avalon_universal_slave_0_agent:m0_address -> key2_s1_translator:uav_address
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // key2_s1_translator_avalon_universal_slave_0_agent:m0_write -> key2_s1_translator:uav_write
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // key2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key2_s1_translator:uav_lock
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // key2_s1_translator_avalon_universal_slave_0_agent:m0_read -> key2_s1_translator:uav_read
	wire  [31:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // key2_s1_translator:uav_readdata -> key2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // key2_s1_translator:uav_readdatavalid -> key2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // key2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key2_s1_translator:uav_debugaccess
	wire   [3:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // key2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key2_s1_translator:uav_byteenable
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] key2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // key1_s1_translator:uav_waitrequest -> key1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // key1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key1_s1_translator:uav_burstcount
	wire  [31:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // key1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key1_s1_translator:uav_writedata
	wire  [20:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // key1_s1_translator_avalon_universal_slave_0_agent:m0_address -> key1_s1_translator:uav_address
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // key1_s1_translator_avalon_universal_slave_0_agent:m0_write -> key1_s1_translator:uav_write
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // key1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key1_s1_translator:uav_lock
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // key1_s1_translator_avalon_universal_slave_0_agent:m0_read -> key1_s1_translator:uav_read
	wire  [31:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // key1_s1_translator:uav_readdata -> key1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // key1_s1_translator:uav_readdatavalid -> key1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // key1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key1_s1_translator:uav_debugaccess
	wire   [3:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // key1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key1_s1_translator:uav_byteenable
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] key1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [20:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // ledr_s1_translator:uav_waitrequest -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // ledr_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ledr_s1_translator:uav_burstcount
	wire  [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // ledr_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ledr_s1_translator:uav_writedata
	wire  [20:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // ledr_s1_translator_avalon_universal_slave_0_agent:m0_address -> ledr_s1_translator:uav_address
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // ledr_s1_translator_avalon_universal_slave_0_agent:m0_write -> ledr_s1_translator:uav_write
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // ledr_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ledr_s1_translator:uav_lock
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // ledr_s1_translator_avalon_universal_slave_0_agent:m0_read -> ledr_s1_translator:uav_read
	wire  [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // ledr_s1_translator:uav_readdata -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // ledr_s1_translator:uav_readdatavalid -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // ledr_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ledr_s1_translator:uav_debugaccess
	wire   [3:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // ledr_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ledr_s1_translator:uav_byteenable
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // LCD_DATA_s1_translator:uav_waitrequest -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_DATA_s1_translator:uav_burstcount
	wire  [31:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_DATA_s1_translator:uav_writedata
	wire  [20:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_address -> LCD_DATA_s1_translator:uav_address
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_write -> LCD_DATA_s1_translator:uav_write
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_DATA_s1_translator:uav_lock
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_read -> LCD_DATA_s1_translator:uav_read
	wire  [31:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // LCD_DATA_s1_translator:uav_readdata -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // LCD_DATA_s1_translator:uav_readdatavalid -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_DATA_s1_translator:uav_debugaccess
	wire   [3:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_DATA_s1_translator:uav_byteenable
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // LCD_RW_s1_translator:uav_waitrequest -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_RW_s1_translator:uav_burstcount
	wire  [31:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_RW_s1_translator:uav_writedata
	wire  [20:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_address -> LCD_RW_s1_translator:uav_address
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_write -> LCD_RW_s1_translator:uav_write
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_RW_s1_translator:uav_lock
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_read -> LCD_RW_s1_translator:uav_read
	wire  [31:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // LCD_RW_s1_translator:uav_readdata -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // LCD_RW_s1_translator:uav_readdatavalid -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_RW_s1_translator:uav_debugaccess
	wire   [3:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // LCD_RW_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_RW_s1_translator:uav_byteenable
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // LCD_RS_s1_translator:uav_waitrequest -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_RS_s1_translator:uav_burstcount
	wire  [31:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_RS_s1_translator:uav_writedata
	wire  [20:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_address -> LCD_RS_s1_translator:uav_address
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_write -> LCD_RS_s1_translator:uav_write
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_RS_s1_translator:uav_lock
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_read -> LCD_RS_s1_translator:uav_read
	wire  [31:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // LCD_RS_s1_translator:uav_readdata -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // LCD_RS_s1_translator:uav_readdatavalid -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_RS_s1_translator:uav_debugaccess
	wire   [3:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // LCD_RS_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_RS_s1_translator:uav_byteenable
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // LCD_EN_s1_translator:uav_waitrequest -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_EN_s1_translator:uav_burstcount
	wire  [31:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_EN_s1_translator:uav_writedata
	wire  [20:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_address -> LCD_EN_s1_translator:uav_address
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_write -> LCD_EN_s1_translator:uav_write
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_EN_s1_translator:uav_lock
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_read -> LCD_EN_s1_translator:uav_read
	wire  [31:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // LCD_EN_s1_translator:uav_readdata -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // LCD_EN_s1_translator:uav_readdatavalid -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_EN_s1_translator:uav_debugaccess
	wire   [3:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // LCD_EN_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_EN_s1_translator:uav_byteenable
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // LCD_ON_s1_translator:uav_waitrequest -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_ON_s1_translator:uav_burstcount
	wire  [31:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_ON_s1_translator:uav_writedata
	wire  [20:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_address -> LCD_ON_s1_translator:uav_address
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_write -> LCD_ON_s1_translator:uav_write
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_ON_s1_translator:uav_lock
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_read -> LCD_ON_s1_translator:uav_read
	wire  [31:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // LCD_ON_s1_translator:uav_readdata -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // LCD_ON_s1_translator:uav_readdatavalid -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_ON_s1_translator:uav_debugaccess
	wire   [3:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // LCD_ON_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_ON_s1_translator:uav_byteenable
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [97:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [97:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [97:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [97:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [97:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_002:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led8_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led8_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led8_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [97:0] led8_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led8_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         led8_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_003:sink_ready -> led8_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led7_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led7_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led7_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [97:0] led7_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led7_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         led7_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_004:sink_ready -> led7_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led6_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led6_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led6_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [97:0] led6_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led6_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         led6_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_005:sink_ready -> led6_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [97:0] led5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         led5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_006:sink_ready -> led5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [97:0] led4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         led4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_007:sink_ready -> led4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [97:0] led3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         led3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_008:sink_ready -> led3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [97:0] led2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         led2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_009:sink_ready -> led2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [97:0] led1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         led1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_010:sink_ready -> led1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [97:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_011:sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // switch0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // switch0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // switch0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [97:0] switch0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // switch0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_012:sink_ready -> switch0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // key3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // key3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // key3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [97:0] key3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // key3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_013:sink_ready -> key3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // key2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // key2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // key2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [97:0] key2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // key2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_014:sink_ready -> key2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // key1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // key1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // key1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [97:0] key1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // key1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_015:sink_ready -> key1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [97:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_016:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // ledr_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // ledr_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // ledr_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [97:0] ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // ledr_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_017:sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [97:0] lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire         lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_018:sink_ready -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [97:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // LCD_RW_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_019:sink_ready -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [97:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // LCD_RS_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_020:sink_ready -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [97:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // LCD_EN_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_021:sink_ready -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [97:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // LCD_ON_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_022:sink_ready -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led1:reset_n, led1_s1_translator:reset, led1_s1_translator_avalon_universal_slave_0_agent:reset, led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led2:reset_n, led2_s1_translator:reset, led2_s1_translator_avalon_universal_slave_0_agent:reset, led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led3:reset_n, led3_s1_translator:reset, led3_s1_translator_avalon_universal_slave_0_agent:reset, led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led4:reset_n, led4_s1_translator:reset, led4_s1_translator_avalon_universal_slave_0_agent:reset, led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led5:reset_n, led5_s1_translator:reset, led5_s1_translator_avalon_universal_slave_0_agent:reset, led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led6:reset_n, led6_s1_translator:reset, led6_s1_translator_avalon_universal_slave_0_agent:reset, led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led7:reset_n, led7_s1_translator:reset, led7_s1_translator_avalon_universal_slave_0_agent:reset, led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led8:reset_n, led8_s1_translator:reset, led8_s1_translator_avalon_universal_slave_0_agent:reset, led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset]
	wire         rst_controller_reset_out_reset_req;                                                                  // rst_controller:reset_req -> onchip_memory2_0:reset_req
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                                          // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                                                  // rst_controller_001:reset_out -> [LCD_DATA:reset_n, LCD_DATA_s1_translator:reset, LCD_DATA_s1_translator_avalon_universal_slave_0_agent:reset, LCD_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_EN:reset_n, LCD_EN_s1_translator:reset, LCD_EN_s1_translator_avalon_universal_slave_0_agent:reset, LCD_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_ON:reset_n, LCD_ON_s1_translator:reset, LCD_ON_s1_translator_avalon_universal_slave_0_agent:reset, LCD_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_RS:reset_n, LCD_RS_s1_translator:reset, LCD_RS_s1_translator_avalon_universal_slave_0_agent:reset, LCD_RS_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_RW:reset_n, LCD_RW_s1_translator:reset, LCD_RW_s1_translator_avalon_universal_slave_0_agent:reset, LCD_RW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_011:reset, cmd_xbar_mux_012:reset, cmd_xbar_mux_013:reset, cmd_xbar_mux_014:reset, cmd_xbar_mux_015:reset, cmd_xbar_mux_016:reset, cmd_xbar_mux_017:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, key1:reset_n, key1_s1_translator:reset, key1_s1_translator_avalon_universal_slave_0_agent:reset, key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key2:reset_n, key2_s1_translator:reset, key2_s1_translator_avalon_universal_slave_0_agent:reset, key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key3:reset_n, key3_s1_translator:reset, key3_s1_translator_avalon_universal_slave_0_agent:reset, key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ledr:reset_n, ledr_s1_translator:reset, ledr_s1_translator_avalon_universal_slave_0_agent:reset, ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, switch0:reset_n, switch0_s1_translator:reset, switch0_s1_translator_avalon_universal_slave_0_agent:reset, switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart_0:reset_n, uart_0_s1_translator:reset, uart_0_s1_translator_avalon_universal_slave_0_agent:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [22:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [22:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                     // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                           // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                   // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src2_data;                                                                            // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [22:0] cmd_xbar_demux_src2_channel;                                                                         // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                           // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                     // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                           // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                   // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src3_data;                                                                            // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire  [22:0] cmd_xbar_demux_src3_channel;                                                                         // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                           // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                     // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                           // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                   // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src4_data;                                                                            // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire  [22:0] cmd_xbar_demux_src4_channel;                                                                         // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                           // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_src5_endofpacket;                                                                     // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                           // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                                   // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src5_data;                                                                            // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire  [22:0] cmd_xbar_demux_src5_channel;                                                                         // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire         cmd_xbar_demux_src5_ready;                                                                           // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire         cmd_xbar_demux_src6_endofpacket;                                                                     // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                           // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                                   // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src6_data;                                                                            // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire  [22:0] cmd_xbar_demux_src6_channel;                                                                         // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire         cmd_xbar_demux_src6_ready;                                                                           // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire         cmd_xbar_demux_src7_endofpacket;                                                                     // cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire         cmd_xbar_demux_src7_valid;                                                                           // cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire         cmd_xbar_demux_src7_startofpacket;                                                                   // cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src7_data;                                                                            // cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	wire  [22:0] cmd_xbar_demux_src7_channel;                                                                         // cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire         cmd_xbar_demux_src7_ready;                                                                           // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire         cmd_xbar_demux_src8_endofpacket;                                                                     // cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire         cmd_xbar_demux_src8_valid;                                                                           // cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire         cmd_xbar_demux_src8_startofpacket;                                                                   // cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src8_data;                                                                            // cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	wire  [22:0] cmd_xbar_demux_src8_channel;                                                                         // cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire         cmd_xbar_demux_src8_ready;                                                                           // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire         cmd_xbar_demux_src9_endofpacket;                                                                     // cmd_xbar_demux:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire         cmd_xbar_demux_src9_valid;                                                                           // cmd_xbar_demux:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire         cmd_xbar_demux_src9_startofpacket;                                                                   // cmd_xbar_demux:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src9_data;                                                                            // cmd_xbar_demux:src9_data -> cmd_xbar_mux_009:sink0_data
	wire  [22:0] cmd_xbar_demux_src9_channel;                                                                         // cmd_xbar_demux:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire         cmd_xbar_demux_src9_ready;                                                                           // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux:src9_ready
	wire         cmd_xbar_demux_src10_endofpacket;                                                                    // cmd_xbar_demux:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire         cmd_xbar_demux_src10_valid;                                                                          // cmd_xbar_demux:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire         cmd_xbar_demux_src10_startofpacket;                                                                  // cmd_xbar_demux:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src10_data;                                                                           // cmd_xbar_demux:src10_data -> cmd_xbar_mux_010:sink0_data
	wire  [22:0] cmd_xbar_demux_src10_channel;                                                                        // cmd_xbar_demux:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire         cmd_xbar_demux_src10_ready;                                                                          // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux:src10_ready
	wire         cmd_xbar_demux_src11_endofpacket;                                                                    // cmd_xbar_demux:src11_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	wire         cmd_xbar_demux_src11_valid;                                                                          // cmd_xbar_demux:src11_valid -> cmd_xbar_mux_011:sink0_valid
	wire         cmd_xbar_demux_src11_startofpacket;                                                                  // cmd_xbar_demux:src11_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src11_data;                                                                           // cmd_xbar_demux:src11_data -> cmd_xbar_mux_011:sink0_data
	wire  [22:0] cmd_xbar_demux_src11_channel;                                                                        // cmd_xbar_demux:src11_channel -> cmd_xbar_mux_011:sink0_channel
	wire         cmd_xbar_demux_src11_ready;                                                                          // cmd_xbar_mux_011:sink0_ready -> cmd_xbar_demux:src11_ready
	wire         cmd_xbar_demux_src12_endofpacket;                                                                    // cmd_xbar_demux:src12_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	wire         cmd_xbar_demux_src12_valid;                                                                          // cmd_xbar_demux:src12_valid -> cmd_xbar_mux_012:sink0_valid
	wire         cmd_xbar_demux_src12_startofpacket;                                                                  // cmd_xbar_demux:src12_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src12_data;                                                                           // cmd_xbar_demux:src12_data -> cmd_xbar_mux_012:sink0_data
	wire  [22:0] cmd_xbar_demux_src12_channel;                                                                        // cmd_xbar_demux:src12_channel -> cmd_xbar_mux_012:sink0_channel
	wire         cmd_xbar_demux_src12_ready;                                                                          // cmd_xbar_mux_012:sink0_ready -> cmd_xbar_demux:src12_ready
	wire         cmd_xbar_demux_src13_endofpacket;                                                                    // cmd_xbar_demux:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire         cmd_xbar_demux_src13_valid;                                                                          // cmd_xbar_demux:src13_valid -> cmd_xbar_mux_013:sink0_valid
	wire         cmd_xbar_demux_src13_startofpacket;                                                                  // cmd_xbar_demux:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src13_data;                                                                           // cmd_xbar_demux:src13_data -> cmd_xbar_mux_013:sink0_data
	wire  [22:0] cmd_xbar_demux_src13_channel;                                                                        // cmd_xbar_demux:src13_channel -> cmd_xbar_mux_013:sink0_channel
	wire         cmd_xbar_demux_src13_ready;                                                                          // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux:src13_ready
	wire         cmd_xbar_demux_src14_endofpacket;                                                                    // cmd_xbar_demux:src14_endofpacket -> cmd_xbar_mux_014:sink0_endofpacket
	wire         cmd_xbar_demux_src14_valid;                                                                          // cmd_xbar_demux:src14_valid -> cmd_xbar_mux_014:sink0_valid
	wire         cmd_xbar_demux_src14_startofpacket;                                                                  // cmd_xbar_demux:src14_startofpacket -> cmd_xbar_mux_014:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src14_data;                                                                           // cmd_xbar_demux:src14_data -> cmd_xbar_mux_014:sink0_data
	wire  [22:0] cmd_xbar_demux_src14_channel;                                                                        // cmd_xbar_demux:src14_channel -> cmd_xbar_mux_014:sink0_channel
	wire         cmd_xbar_demux_src14_ready;                                                                          // cmd_xbar_mux_014:sink0_ready -> cmd_xbar_demux:src14_ready
	wire         cmd_xbar_demux_src15_endofpacket;                                                                    // cmd_xbar_demux:src15_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	wire         cmd_xbar_demux_src15_valid;                                                                          // cmd_xbar_demux:src15_valid -> cmd_xbar_mux_015:sink0_valid
	wire         cmd_xbar_demux_src15_startofpacket;                                                                  // cmd_xbar_demux:src15_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src15_data;                                                                           // cmd_xbar_demux:src15_data -> cmd_xbar_mux_015:sink0_data
	wire  [22:0] cmd_xbar_demux_src15_channel;                                                                        // cmd_xbar_demux:src15_channel -> cmd_xbar_mux_015:sink0_channel
	wire         cmd_xbar_demux_src15_ready;                                                                          // cmd_xbar_mux_015:sink0_ready -> cmd_xbar_demux:src15_ready
	wire         cmd_xbar_demux_src16_endofpacket;                                                                    // cmd_xbar_demux:src16_endofpacket -> cmd_xbar_mux_016:sink0_endofpacket
	wire         cmd_xbar_demux_src16_valid;                                                                          // cmd_xbar_demux:src16_valid -> cmd_xbar_mux_016:sink0_valid
	wire         cmd_xbar_demux_src16_startofpacket;                                                                  // cmd_xbar_demux:src16_startofpacket -> cmd_xbar_mux_016:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src16_data;                                                                           // cmd_xbar_demux:src16_data -> cmd_xbar_mux_016:sink0_data
	wire  [22:0] cmd_xbar_demux_src16_channel;                                                                        // cmd_xbar_demux:src16_channel -> cmd_xbar_mux_016:sink0_channel
	wire         cmd_xbar_demux_src16_ready;                                                                          // cmd_xbar_mux_016:sink0_ready -> cmd_xbar_demux:src16_ready
	wire         cmd_xbar_demux_src17_endofpacket;                                                                    // cmd_xbar_demux:src17_endofpacket -> cmd_xbar_mux_017:sink0_endofpacket
	wire         cmd_xbar_demux_src17_valid;                                                                          // cmd_xbar_demux:src17_valid -> cmd_xbar_mux_017:sink0_valid
	wire         cmd_xbar_demux_src17_startofpacket;                                                                  // cmd_xbar_demux:src17_startofpacket -> cmd_xbar_mux_017:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src17_data;                                                                           // cmd_xbar_demux:src17_data -> cmd_xbar_mux_017:sink0_data
	wire  [22:0] cmd_xbar_demux_src17_channel;                                                                        // cmd_xbar_demux:src17_channel -> cmd_xbar_mux_017:sink0_channel
	wire         cmd_xbar_demux_src17_ready;                                                                          // cmd_xbar_mux_017:sink0_ready -> cmd_xbar_demux:src17_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                       // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                 // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                       // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                               // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src3_data;                                                                        // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src3_channel;                                                                     // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                       // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                 // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                       // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                               // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src4_data;                                                                        // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src4_channel;                                                                     // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                       // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                 // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                       // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                               // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src5_data;                                                                        // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src5_channel;                                                                     // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                       // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                 // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                       // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                               // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src6_data;                                                                        // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src6_channel;                                                                     // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                       // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                 // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                       // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                               // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src7_data;                                                                        // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src7_channel;                                                                     // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	wire         cmd_xbar_demux_001_src7_ready;                                                                       // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                 // cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                       // cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink1_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                               // cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src8_data;                                                                        // cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src8_channel;                                                                     // cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink1_channel
	wire         cmd_xbar_demux_001_src8_ready;                                                                       // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src8_ready
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                 // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                       // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink1_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                               // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src9_data;                                                                        // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src9_channel;                                                                     // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink1_channel
	wire         cmd_xbar_demux_001_src9_ready;                                                                       // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_001:src9_ready
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                      // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink1_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                              // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src10_data;                                                                       // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src10_channel;                                                                    // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink1_channel
	wire         cmd_xbar_demux_001_src10_ready;                                                                      // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_001:src10_ready
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                                // cmd_xbar_demux_001:src11_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                      // cmd_xbar_demux_001:src11_valid -> cmd_xbar_mux_011:sink1_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                              // cmd_xbar_demux_001:src11_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src11_data;                                                                       // cmd_xbar_demux_001:src11_data -> cmd_xbar_mux_011:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src11_channel;                                                                    // cmd_xbar_demux_001:src11_channel -> cmd_xbar_mux_011:sink1_channel
	wire         cmd_xbar_demux_001_src11_ready;                                                                      // cmd_xbar_mux_011:sink1_ready -> cmd_xbar_demux_001:src11_ready
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                                // cmd_xbar_demux_001:src12_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                      // cmd_xbar_demux_001:src12_valid -> cmd_xbar_mux_012:sink1_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                              // cmd_xbar_demux_001:src12_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src12_data;                                                                       // cmd_xbar_demux_001:src12_data -> cmd_xbar_mux_012:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src12_channel;                                                                    // cmd_xbar_demux_001:src12_channel -> cmd_xbar_mux_012:sink1_channel
	wire         cmd_xbar_demux_001_src12_ready;                                                                      // cmd_xbar_mux_012:sink1_ready -> cmd_xbar_demux_001:src12_ready
	wire         cmd_xbar_demux_001_src13_endofpacket;                                                                // cmd_xbar_demux_001:src13_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire         cmd_xbar_demux_001_src13_valid;                                                                      // cmd_xbar_demux_001:src13_valid -> cmd_xbar_mux_013:sink1_valid
	wire         cmd_xbar_demux_001_src13_startofpacket;                                                              // cmd_xbar_demux_001:src13_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src13_data;                                                                       // cmd_xbar_demux_001:src13_data -> cmd_xbar_mux_013:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src13_channel;                                                                    // cmd_xbar_demux_001:src13_channel -> cmd_xbar_mux_013:sink1_channel
	wire         cmd_xbar_demux_001_src13_ready;                                                                      // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_001:src13_ready
	wire         cmd_xbar_demux_001_src14_endofpacket;                                                                // cmd_xbar_demux_001:src14_endofpacket -> cmd_xbar_mux_014:sink1_endofpacket
	wire         cmd_xbar_demux_001_src14_valid;                                                                      // cmd_xbar_demux_001:src14_valid -> cmd_xbar_mux_014:sink1_valid
	wire         cmd_xbar_demux_001_src14_startofpacket;                                                              // cmd_xbar_demux_001:src14_startofpacket -> cmd_xbar_mux_014:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src14_data;                                                                       // cmd_xbar_demux_001:src14_data -> cmd_xbar_mux_014:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src14_channel;                                                                    // cmd_xbar_demux_001:src14_channel -> cmd_xbar_mux_014:sink1_channel
	wire         cmd_xbar_demux_001_src14_ready;                                                                      // cmd_xbar_mux_014:sink1_ready -> cmd_xbar_demux_001:src14_ready
	wire         cmd_xbar_demux_001_src15_endofpacket;                                                                // cmd_xbar_demux_001:src15_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	wire         cmd_xbar_demux_001_src15_valid;                                                                      // cmd_xbar_demux_001:src15_valid -> cmd_xbar_mux_015:sink1_valid
	wire         cmd_xbar_demux_001_src15_startofpacket;                                                              // cmd_xbar_demux_001:src15_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src15_data;                                                                       // cmd_xbar_demux_001:src15_data -> cmd_xbar_mux_015:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src15_channel;                                                                    // cmd_xbar_demux_001:src15_channel -> cmd_xbar_mux_015:sink1_channel
	wire         cmd_xbar_demux_001_src15_ready;                                                                      // cmd_xbar_mux_015:sink1_ready -> cmd_xbar_demux_001:src15_ready
	wire         cmd_xbar_demux_001_src16_endofpacket;                                                                // cmd_xbar_demux_001:src16_endofpacket -> cmd_xbar_mux_016:sink1_endofpacket
	wire         cmd_xbar_demux_001_src16_valid;                                                                      // cmd_xbar_demux_001:src16_valid -> cmd_xbar_mux_016:sink1_valid
	wire         cmd_xbar_demux_001_src16_startofpacket;                                                              // cmd_xbar_demux_001:src16_startofpacket -> cmd_xbar_mux_016:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src16_data;                                                                       // cmd_xbar_demux_001:src16_data -> cmd_xbar_mux_016:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src16_channel;                                                                    // cmd_xbar_demux_001:src16_channel -> cmd_xbar_mux_016:sink1_channel
	wire         cmd_xbar_demux_001_src16_ready;                                                                      // cmd_xbar_mux_016:sink1_ready -> cmd_xbar_demux_001:src16_ready
	wire         cmd_xbar_demux_001_src17_endofpacket;                                                                // cmd_xbar_demux_001:src17_endofpacket -> cmd_xbar_mux_017:sink1_endofpacket
	wire         cmd_xbar_demux_001_src17_valid;                                                                      // cmd_xbar_demux_001:src17_valid -> cmd_xbar_mux_017:sink1_valid
	wire         cmd_xbar_demux_001_src17_startofpacket;                                                              // cmd_xbar_demux_001:src17_startofpacket -> cmd_xbar_mux_017:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src17_data;                                                                       // cmd_xbar_demux_001:src17_data -> cmd_xbar_mux_017:sink1_data
	wire  [22:0] cmd_xbar_demux_001_src17_channel;                                                                    // cmd_xbar_demux_001:src17_channel -> cmd_xbar_mux_017:sink1_channel
	wire         cmd_xbar_demux_001_src17_ready;                                                                      // cmd_xbar_mux_017:sink1_ready -> cmd_xbar_demux_001:src17_ready
	wire         cmd_xbar_demux_001_src18_endofpacket;                                                                // cmd_xbar_demux_001:src18_endofpacket -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src18_valid;                                                                      // cmd_xbar_demux_001:src18_valid -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src18_startofpacket;                                                              // cmd_xbar_demux_001:src18_startofpacket -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src18_data;                                                                       // cmd_xbar_demux_001:src18_data -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_demux_001_src18_channel;                                                                    // cmd_xbar_demux_001:src18_channel -> LCD_DATA_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src19_endofpacket;                                                                // cmd_xbar_demux_001:src19_endofpacket -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src19_valid;                                                                      // cmd_xbar_demux_001:src19_valid -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src19_startofpacket;                                                              // cmd_xbar_demux_001:src19_startofpacket -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src19_data;                                                                       // cmd_xbar_demux_001:src19_data -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_demux_001_src19_channel;                                                                    // cmd_xbar_demux_001:src19_channel -> LCD_RW_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src20_endofpacket;                                                                // cmd_xbar_demux_001:src20_endofpacket -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src20_valid;                                                                      // cmd_xbar_demux_001:src20_valid -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src20_startofpacket;                                                              // cmd_xbar_demux_001:src20_startofpacket -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src20_data;                                                                       // cmd_xbar_demux_001:src20_data -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_demux_001_src20_channel;                                                                    // cmd_xbar_demux_001:src20_channel -> LCD_RS_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src21_endofpacket;                                                                // cmd_xbar_demux_001:src21_endofpacket -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src21_valid;                                                                      // cmd_xbar_demux_001:src21_valid -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src21_startofpacket;                                                              // cmd_xbar_demux_001:src21_startofpacket -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src21_data;                                                                       // cmd_xbar_demux_001:src21_data -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_demux_001_src21_channel;                                                                    // cmd_xbar_demux_001:src21_channel -> LCD_EN_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src22_endofpacket;                                                                // cmd_xbar_demux_001:src22_endofpacket -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src22_valid;                                                                      // cmd_xbar_demux_001:src22_valid -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src22_startofpacket;                                                              // cmd_xbar_demux_001:src22_startofpacket -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src22_data;                                                                       // cmd_xbar_demux_001:src22_data -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_demux_001_src22_channel;                                                                    // cmd_xbar_demux_001:src22_channel -> LCD_ON_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [97:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [22:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [97:0] rsp_xbar_demux_src1_data;                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [22:0] rsp_xbar_demux_src1_channel;                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                           // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [97:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [22:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                 // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                       // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                               // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [97:0] rsp_xbar_demux_001_src1_data;                                                                        // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [22:0] rsp_xbar_demux_001_src1_channel;                                                                     // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [97:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [22:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                       // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                 // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                       // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                               // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [97:0] rsp_xbar_demux_002_src1_data;                                                                        // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [22:0] rsp_xbar_demux_002_src1_channel;                                                                     // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [97:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire  [22:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                       // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                 // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                       // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                               // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [97:0] rsp_xbar_demux_003_src1_data;                                                                        // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire  [22:0] rsp_xbar_demux_003_src1_channel;                                                                     // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                       // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [97:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire  [22:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                       // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                 // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                       // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                               // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [97:0] rsp_xbar_demux_004_src1_data;                                                                        // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire  [22:0] rsp_xbar_demux_004_src1_channel;                                                                     // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                       // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [97:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire  [22:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_005_src1_endofpacket;                                                                 // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src1_valid;                                                                       // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src1_startofpacket;                                                               // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [97:0] rsp_xbar_demux_005_src1_data;                                                                        // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire  [22:0] rsp_xbar_demux_005_src1_channel;                                                                     // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src1_ready;                                                                       // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                 // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                       // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                               // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [97:0] rsp_xbar_demux_006_src0_data;                                                                        // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire  [22:0] rsp_xbar_demux_006_src0_channel;                                                                     // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                       // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_006_src1_endofpacket;                                                                 // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src1_valid;                                                                       // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src1_startofpacket;                                                               // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [97:0] rsp_xbar_demux_006_src1_data;                                                                        // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	wire  [22:0] rsp_xbar_demux_006_src1_channel;                                                                     // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src1_ready;                                                                       // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                 // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                       // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                               // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [97:0] rsp_xbar_demux_007_src0_data;                                                                        // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire  [22:0] rsp_xbar_demux_007_src0_channel;                                                                     // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                       // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_007_src1_endofpacket;                                                                 // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src1_valid;                                                                       // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src1_startofpacket;                                                               // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [97:0] rsp_xbar_demux_007_src1_data;                                                                        // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	wire  [22:0] rsp_xbar_demux_007_src1_channel;                                                                     // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src1_ready;                                                                       // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                 // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                       // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                               // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [97:0] rsp_xbar_demux_008_src0_data;                                                                        // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire  [22:0] rsp_xbar_demux_008_src0_channel;                                                                     // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                       // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_008_src1_endofpacket;                                                                 // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src1_valid;                                                                       // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src1_startofpacket;                                                               // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [97:0] rsp_xbar_demux_008_src1_data;                                                                        // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink8_data
	wire  [22:0] rsp_xbar_demux_008_src1_channel;                                                                     // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src1_ready;                                                                       // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src1_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                 // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                       // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                               // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [97:0] rsp_xbar_demux_009_src0_data;                                                                        // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire  [22:0] rsp_xbar_demux_009_src0_channel;                                                                     // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                       // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_009_src1_endofpacket;                                                                 // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src1_valid;                                                                       // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src1_startofpacket;                                                               // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [97:0] rsp_xbar_demux_009_src1_data;                                                                        // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_001:sink9_data
	wire  [22:0] rsp_xbar_demux_009_src1_channel;                                                                     // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src1_ready;                                                                       // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src1_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                 // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                       // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                               // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [97:0] rsp_xbar_demux_010_src0_data;                                                                        // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire  [22:0] rsp_xbar_demux_010_src0_channel;                                                                     // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                       // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_010_src1_endofpacket;                                                                 // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src1_valid;                                                                       // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src1_startofpacket;                                                               // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [97:0] rsp_xbar_demux_010_src1_data;                                                                        // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_001:sink10_data
	wire  [22:0] rsp_xbar_demux_010_src1_channel;                                                                     // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src1_ready;                                                                       // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src1_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                 // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                       // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                               // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	wire  [97:0] rsp_xbar_demux_011_src0_data;                                                                        // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	wire  [22:0] rsp_xbar_demux_011_src0_channel;                                                                     // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                       // rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_011_src1_endofpacket;                                                                 // rsp_xbar_demux_011:src1_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src1_valid;                                                                       // rsp_xbar_demux_011:src1_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src1_startofpacket;                                                               // rsp_xbar_demux_011:src1_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [97:0] rsp_xbar_demux_011_src1_data;                                                                        // rsp_xbar_demux_011:src1_data -> rsp_xbar_mux_001:sink11_data
	wire  [22:0] rsp_xbar_demux_011_src1_channel;                                                                     // rsp_xbar_demux_011:src1_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src1_ready;                                                                       // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src1_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                 // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                       // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                               // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	wire  [97:0] rsp_xbar_demux_012_src0_data;                                                                        // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	wire  [22:0] rsp_xbar_demux_012_src0_channel;                                                                     // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                       // rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_012_src1_endofpacket;                                                                 // rsp_xbar_demux_012:src1_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src1_valid;                                                                       // rsp_xbar_demux_012:src1_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src1_startofpacket;                                                               // rsp_xbar_demux_012:src1_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [97:0] rsp_xbar_demux_012_src1_data;                                                                        // rsp_xbar_demux_012:src1_data -> rsp_xbar_mux_001:sink12_data
	wire  [22:0] rsp_xbar_demux_012_src1_channel;                                                                     // rsp_xbar_demux_012:src1_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src1_ready;                                                                       // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src1_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                 // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                       // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                               // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	wire  [97:0] rsp_xbar_demux_013_src0_data;                                                                        // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	wire  [22:0] rsp_xbar_demux_013_src0_channel;                                                                     // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                       // rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_013_src1_endofpacket;                                                                 // rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire         rsp_xbar_demux_013_src1_valid;                                                                       // rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_001:sink13_valid
	wire         rsp_xbar_demux_013_src1_startofpacket;                                                               // rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [97:0] rsp_xbar_demux_013_src1_data;                                                                        // rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_001:sink13_data
	wire  [22:0] rsp_xbar_demux_013_src1_channel;                                                                     // rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_001:sink13_channel
	wire         rsp_xbar_demux_013_src1_ready;                                                                       // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src1_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                                 // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                       // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                               // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	wire  [97:0] rsp_xbar_demux_014_src0_data;                                                                        // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	wire  [22:0] rsp_xbar_demux_014_src0_channel;                                                                     // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                       // rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_014_src1_endofpacket;                                                                 // rsp_xbar_demux_014:src1_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire         rsp_xbar_demux_014_src1_valid;                                                                       // rsp_xbar_demux_014:src1_valid -> rsp_xbar_mux_001:sink14_valid
	wire         rsp_xbar_demux_014_src1_startofpacket;                                                               // rsp_xbar_demux_014:src1_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [97:0] rsp_xbar_demux_014_src1_data;                                                                        // rsp_xbar_demux_014:src1_data -> rsp_xbar_mux_001:sink14_data
	wire  [22:0] rsp_xbar_demux_014_src1_channel;                                                                     // rsp_xbar_demux_014:src1_channel -> rsp_xbar_mux_001:sink14_channel
	wire         rsp_xbar_demux_014_src1_ready;                                                                       // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src1_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                                 // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                       // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                               // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	wire  [97:0] rsp_xbar_demux_015_src0_data;                                                                        // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux:sink15_data
	wire  [22:0] rsp_xbar_demux_015_src0_channel;                                                                     // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                       // rsp_xbar_mux:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_015_src1_endofpacket;                                                                 // rsp_xbar_demux_015:src1_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire         rsp_xbar_demux_015_src1_valid;                                                                       // rsp_xbar_demux_015:src1_valid -> rsp_xbar_mux_001:sink15_valid
	wire         rsp_xbar_demux_015_src1_startofpacket;                                                               // rsp_xbar_demux_015:src1_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [97:0] rsp_xbar_demux_015_src1_data;                                                                        // rsp_xbar_demux_015:src1_data -> rsp_xbar_mux_001:sink15_data
	wire  [22:0] rsp_xbar_demux_015_src1_channel;                                                                     // rsp_xbar_demux_015:src1_channel -> rsp_xbar_mux_001:sink15_channel
	wire         rsp_xbar_demux_015_src1_ready;                                                                       // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src1_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                                 // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                       // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                               // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux:sink16_startofpacket
	wire  [97:0] rsp_xbar_demux_016_src0_data;                                                                        // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux:sink16_data
	wire  [22:0] rsp_xbar_demux_016_src0_channel;                                                                     // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                       // rsp_xbar_mux:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_016_src1_endofpacket;                                                                 // rsp_xbar_demux_016:src1_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire         rsp_xbar_demux_016_src1_valid;                                                                       // rsp_xbar_demux_016:src1_valid -> rsp_xbar_mux_001:sink16_valid
	wire         rsp_xbar_demux_016_src1_startofpacket;                                                               // rsp_xbar_demux_016:src1_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [97:0] rsp_xbar_demux_016_src1_data;                                                                        // rsp_xbar_demux_016:src1_data -> rsp_xbar_mux_001:sink16_data
	wire  [22:0] rsp_xbar_demux_016_src1_channel;                                                                     // rsp_xbar_demux_016:src1_channel -> rsp_xbar_mux_001:sink16_channel
	wire         rsp_xbar_demux_016_src1_ready;                                                                       // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src1_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                                 // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                                       // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                               // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux:sink17_startofpacket
	wire  [97:0] rsp_xbar_demux_017_src0_data;                                                                        // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux:sink17_data
	wire  [22:0] rsp_xbar_demux_017_src0_channel;                                                                     // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                                       // rsp_xbar_mux:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         rsp_xbar_demux_017_src1_endofpacket;                                                                 // rsp_xbar_demux_017:src1_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire         rsp_xbar_demux_017_src1_valid;                                                                       // rsp_xbar_demux_017:src1_valid -> rsp_xbar_mux_001:sink17_valid
	wire         rsp_xbar_demux_017_src1_startofpacket;                                                               // rsp_xbar_demux_017:src1_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [97:0] rsp_xbar_demux_017_src1_data;                                                                        // rsp_xbar_demux_017:src1_data -> rsp_xbar_mux_001:sink17_data
	wire  [22:0] rsp_xbar_demux_017_src1_channel;                                                                     // rsp_xbar_demux_017:src1_channel -> rsp_xbar_mux_001:sink17_channel
	wire         rsp_xbar_demux_017_src1_ready;                                                                       // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src1_ready
	wire         rsp_xbar_demux_018_src0_endofpacket;                                                                 // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire         rsp_xbar_demux_018_src0_valid;                                                                       // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire         rsp_xbar_demux_018_src0_startofpacket;                                                               // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [97:0] rsp_xbar_demux_018_src0_data;                                                                        // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire  [22:0] rsp_xbar_demux_018_src0_channel;                                                                     // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire         rsp_xbar_demux_018_src0_ready;                                                                       // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire         rsp_xbar_demux_019_src0_endofpacket;                                                                 // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire         rsp_xbar_demux_019_src0_valid;                                                                       // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire         rsp_xbar_demux_019_src0_startofpacket;                                                               // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [97:0] rsp_xbar_demux_019_src0_data;                                                                        // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire  [22:0] rsp_xbar_demux_019_src0_channel;                                                                     // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire         rsp_xbar_demux_019_src0_ready;                                                                       // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire         rsp_xbar_demux_020_src0_endofpacket;                                                                 // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire         rsp_xbar_demux_020_src0_valid;                                                                       // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire         rsp_xbar_demux_020_src0_startofpacket;                                                               // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [97:0] rsp_xbar_demux_020_src0_data;                                                                        // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire  [22:0] rsp_xbar_demux_020_src0_channel;                                                                     // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire         rsp_xbar_demux_020_src0_ready;                                                                       // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire         rsp_xbar_demux_021_src0_endofpacket;                                                                 // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire         rsp_xbar_demux_021_src0_valid;                                                                       // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire         rsp_xbar_demux_021_src0_startofpacket;                                                               // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [97:0] rsp_xbar_demux_021_src0_data;                                                                        // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire  [22:0] rsp_xbar_demux_021_src0_channel;                                                                     // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire         rsp_xbar_demux_021_src0_ready;                                                                       // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire         rsp_xbar_demux_022_src0_endofpacket;                                                                 // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire         rsp_xbar_demux_022_src0_valid;                                                                       // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	wire         rsp_xbar_demux_022_src0_startofpacket;                                                               // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [97:0] rsp_xbar_demux_022_src0_data;                                                                        // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	wire  [22:0] rsp_xbar_demux_022_src0_channel;                                                                     // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	wire         rsp_xbar_demux_022_src0_ready;                                                                       // rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire         addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                               // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [97:0] addr_router_src_data;                                                                                // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire  [22:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [97:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [22:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                              // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [97:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire  [22:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [97:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [22:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                          // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                        // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                              // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                      // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_src_data;                                                                               // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_src_channel;                                                                            // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [97:0] id_router_src_data;                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [22:0] id_router_src_channel;                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                    // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                          // cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                  // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_001_src_data;                                                                           // cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_001_src_channel;                                                                        // cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                             // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [97:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [22:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                             // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                    // cmd_xbar_mux_002:src_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                          // cmd_xbar_mux_002:src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                  // cmd_xbar_mux_002:src_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_002_src_data;                                                                           // cmd_xbar_mux_002:src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_002_src_channel;                                                                        // cmd_xbar_mux_002:src_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [97:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [22:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                    // cmd_xbar_mux_003:src_endofpacket -> led8_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                          // cmd_xbar_mux_003:src_valid -> led8_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                  // cmd_xbar_mux_003:src_startofpacket -> led8_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_003_src_data;                                                                           // cmd_xbar_mux_003:src_data -> led8_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_003_src_channel;                                                                        // cmd_xbar_mux_003:src_channel -> led8_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                          // led8_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [97:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [22:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                    // cmd_xbar_mux_004:src_endofpacket -> led7_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                          // cmd_xbar_mux_004:src_valid -> led7_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                  // cmd_xbar_mux_004:src_startofpacket -> led7_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_004_src_data;                                                                           // cmd_xbar_mux_004:src_data -> led7_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_004_src_channel;                                                                        // cmd_xbar_mux_004:src_channel -> led7_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                          // led7_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire         id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [97:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [22:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_mux_005_src_endofpacket;                                                                    // cmd_xbar_mux_005:src_endofpacket -> led6_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_005_src_valid;                                                                          // cmd_xbar_mux_005:src_valid -> led6_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_005_src_startofpacket;                                                                  // cmd_xbar_mux_005:src_startofpacket -> led6_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_005_src_data;                                                                           // cmd_xbar_mux_005:src_data -> led6_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_005_src_channel;                                                                        // cmd_xbar_mux_005:src_channel -> led6_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_005_src_ready;                                                                          // led6_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire         id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [97:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [22:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_mux_006_src_endofpacket;                                                                    // cmd_xbar_mux_006:src_endofpacket -> led5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_006_src_valid;                                                                          // cmd_xbar_mux_006:src_valid -> led5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_006_src_startofpacket;                                                                  // cmd_xbar_mux_006:src_startofpacket -> led5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_006_src_data;                                                                           // cmd_xbar_mux_006:src_data -> led5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_006_src_channel;                                                                        // cmd_xbar_mux_006:src_channel -> led5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_006_src_ready;                                                                          // led5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire         id_router_006_src_endofpacket;                                                                       // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                             // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                     // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [97:0] id_router_006_src_data;                                                                              // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [22:0] id_router_006_src_channel;                                                                           // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                             // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_007_src_endofpacket;                                                                    // cmd_xbar_mux_007:src_endofpacket -> led4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_007_src_valid;                                                                          // cmd_xbar_mux_007:src_valid -> led4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_007_src_startofpacket;                                                                  // cmd_xbar_mux_007:src_startofpacket -> led4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_007_src_data;                                                                           // cmd_xbar_mux_007:src_data -> led4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_007_src_channel;                                                                        // cmd_xbar_mux_007:src_channel -> led4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_007_src_ready;                                                                          // led4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire         id_router_007_src_endofpacket;                                                                       // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                             // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                     // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [97:0] id_router_007_src_data;                                                                              // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [22:0] id_router_007_src_channel;                                                                           // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                             // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_mux_008_src_endofpacket;                                                                    // cmd_xbar_mux_008:src_endofpacket -> led3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_008_src_valid;                                                                          // cmd_xbar_mux_008:src_valid -> led3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_008_src_startofpacket;                                                                  // cmd_xbar_mux_008:src_startofpacket -> led3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_008_src_data;                                                                           // cmd_xbar_mux_008:src_data -> led3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_008_src_channel;                                                                        // cmd_xbar_mux_008:src_channel -> led3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_008_src_ready;                                                                          // led3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire         id_router_008_src_endofpacket;                                                                       // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                             // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                     // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [97:0] id_router_008_src_data;                                                                              // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [22:0] id_router_008_src_channel;                                                                           // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                             // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_mux_009_src_endofpacket;                                                                    // cmd_xbar_mux_009:src_endofpacket -> led2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_009_src_valid;                                                                          // cmd_xbar_mux_009:src_valid -> led2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_009_src_startofpacket;                                                                  // cmd_xbar_mux_009:src_startofpacket -> led2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_009_src_data;                                                                           // cmd_xbar_mux_009:src_data -> led2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_009_src_channel;                                                                        // cmd_xbar_mux_009:src_channel -> led2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_009_src_ready;                                                                          // led2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire         id_router_009_src_endofpacket;                                                                       // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                             // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                     // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [97:0] id_router_009_src_data;                                                                              // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [22:0] id_router_009_src_channel;                                                                           // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                             // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_mux_010_src_endofpacket;                                                                    // cmd_xbar_mux_010:src_endofpacket -> led1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_010_src_valid;                                                                          // cmd_xbar_mux_010:src_valid -> led1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_010_src_startofpacket;                                                                  // cmd_xbar_mux_010:src_startofpacket -> led1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_010_src_data;                                                                           // cmd_xbar_mux_010:src_data -> led1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_010_src_channel;                                                                        // cmd_xbar_mux_010:src_channel -> led1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_010_src_ready;                                                                          // led1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire         id_router_010_src_endofpacket;                                                                       // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                             // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                     // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [97:0] id_router_010_src_data;                                                                              // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [22:0] id_router_010_src_channel;                                                                           // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                             // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_mux_011_src_endofpacket;                                                                    // cmd_xbar_mux_011:src_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_011_src_valid;                                                                          // cmd_xbar_mux_011:src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_011_src_startofpacket;                                                                  // cmd_xbar_mux_011:src_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_011_src_data;                                                                           // cmd_xbar_mux_011:src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_011_src_channel;                                                                        // cmd_xbar_mux_011:src_channel -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_011_src_ready;                                                                          // uart_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_011:src_ready
	wire         id_router_011_src_endofpacket;                                                                       // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                             // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                     // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [97:0] id_router_011_src_data;                                                                              // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [22:0] id_router_011_src_channel;                                                                           // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                             // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_mux_012_src_endofpacket;                                                                    // cmd_xbar_mux_012:src_endofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_012_src_valid;                                                                          // cmd_xbar_mux_012:src_valid -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_012_src_startofpacket;                                                                  // cmd_xbar_mux_012:src_startofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_012_src_data;                                                                           // cmd_xbar_mux_012:src_data -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_012_src_channel;                                                                        // cmd_xbar_mux_012:src_channel -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_012_src_ready;                                                                          // switch0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_012:src_ready
	wire         id_router_012_src_endofpacket;                                                                       // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                             // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                     // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [97:0] id_router_012_src_data;                                                                              // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [22:0] id_router_012_src_channel;                                                                           // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                             // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_mux_013_src_endofpacket;                                                                    // cmd_xbar_mux_013:src_endofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_013_src_valid;                                                                          // cmd_xbar_mux_013:src_valid -> key3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_013_src_startofpacket;                                                                  // cmd_xbar_mux_013:src_startofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_013_src_data;                                                                           // cmd_xbar_mux_013:src_data -> key3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_013_src_channel;                                                                        // cmd_xbar_mux_013:src_channel -> key3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_013_src_ready;                                                                          // key3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire         id_router_013_src_endofpacket;                                                                       // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                             // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                     // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [97:0] id_router_013_src_data;                                                                              // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [22:0] id_router_013_src_channel;                                                                           // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                             // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_mux_014_src_endofpacket;                                                                    // cmd_xbar_mux_014:src_endofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_014_src_valid;                                                                          // cmd_xbar_mux_014:src_valid -> key2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_014_src_startofpacket;                                                                  // cmd_xbar_mux_014:src_startofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_014_src_data;                                                                           // cmd_xbar_mux_014:src_data -> key2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_014_src_channel;                                                                        // cmd_xbar_mux_014:src_channel -> key2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_014_src_ready;                                                                          // key2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_014:src_ready
	wire         id_router_014_src_endofpacket;                                                                       // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                             // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                     // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [97:0] id_router_014_src_data;                                                                              // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire  [22:0] id_router_014_src_channel;                                                                           // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                             // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_mux_015_src_endofpacket;                                                                    // cmd_xbar_mux_015:src_endofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_015_src_valid;                                                                          // cmd_xbar_mux_015:src_valid -> key1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_015_src_startofpacket;                                                                  // cmd_xbar_mux_015:src_startofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_015_src_data;                                                                           // cmd_xbar_mux_015:src_data -> key1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_015_src_channel;                                                                        // cmd_xbar_mux_015:src_channel -> key1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_015_src_ready;                                                                          // key1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_015:src_ready
	wire         id_router_015_src_endofpacket;                                                                       // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                             // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                     // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [97:0] id_router_015_src_data;                                                                              // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire  [22:0] id_router_015_src_channel;                                                                           // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                             // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_mux_016_src_endofpacket;                                                                    // cmd_xbar_mux_016:src_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_016_src_valid;                                                                          // cmd_xbar_mux_016:src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_016_src_startofpacket;                                                                  // cmd_xbar_mux_016:src_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_016_src_data;                                                                           // cmd_xbar_mux_016:src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_016_src_channel;                                                                        // cmd_xbar_mux_016:src_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_016_src_ready;                                                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_016:src_ready
	wire         id_router_016_src_endofpacket;                                                                       // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                             // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                     // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [97:0] id_router_016_src_data;                                                                              // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire  [22:0] id_router_016_src_channel;                                                                           // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                             // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_mux_017_src_endofpacket;                                                                    // cmd_xbar_mux_017:src_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_017_src_valid;                                                                          // cmd_xbar_mux_017:src_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_017_src_startofpacket;                                                                  // cmd_xbar_mux_017:src_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_017_src_data;                                                                           // cmd_xbar_mux_017:src_data -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [22:0] cmd_xbar_mux_017_src_channel;                                                                        // cmd_xbar_mux_017:src_channel -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_017_src_ready;                                                                          // ledr_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_017:src_ready
	wire         id_router_017_src_endofpacket;                                                                       // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         id_router_017_src_valid;                                                                             // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire         id_router_017_src_startofpacket;                                                                     // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [97:0] id_router_017_src_data;                                                                              // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire  [22:0] id_router_017_src_channel;                                                                           // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire         id_router_017_src_ready;                                                                             // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire         cmd_xbar_demux_001_src18_ready;                                                                      // LCD_DATA_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire         id_router_018_src_endofpacket;                                                                       // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire         id_router_018_src_valid;                                                                             // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire         id_router_018_src_startofpacket;                                                                     // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [97:0] id_router_018_src_data;                                                                              // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire  [22:0] id_router_018_src_channel;                                                                           // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire         id_router_018_src_ready;                                                                             // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire         cmd_xbar_demux_001_src19_ready;                                                                      // LCD_RW_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire         id_router_019_src_endofpacket;                                                                       // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire         id_router_019_src_valid;                                                                             // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire         id_router_019_src_startofpacket;                                                                     // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [97:0] id_router_019_src_data;                                                                              // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire  [22:0] id_router_019_src_channel;                                                                           // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire         id_router_019_src_ready;                                                                             // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire         cmd_xbar_demux_001_src20_ready;                                                                      // LCD_RS_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	wire         id_router_020_src_endofpacket;                                                                       // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire         id_router_020_src_valid;                                                                             // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire         id_router_020_src_startofpacket;                                                                     // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [97:0] id_router_020_src_data;                                                                              // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire  [22:0] id_router_020_src_channel;                                                                           // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire         id_router_020_src_ready;                                                                             // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire         cmd_xbar_demux_001_src21_ready;                                                                      // LCD_EN_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	wire         id_router_021_src_endofpacket;                                                                       // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire         id_router_021_src_valid;                                                                             // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire         id_router_021_src_startofpacket;                                                                     // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [97:0] id_router_021_src_data;                                                                              // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire  [22:0] id_router_021_src_channel;                                                                           // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire         id_router_021_src_ready;                                                                             // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire         cmd_xbar_demux_001_src22_ready;                                                                      // LCD_ON_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	wire         id_router_022_src_endofpacket;                                                                       // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire         id_router_022_src_valid;                                                                             // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire         id_router_022_src_startofpacket;                                                                     // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [97:0] id_router_022_src_data;                                                                              // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire  [22:0] id_router_022_src_channel;                                                                           // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire         id_router_022_src_ready;                                                                             // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire         irq_mapper_receiver0_irq;                                                                            // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                            // uart_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                            // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                            // switch0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	nios_sys_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                                   //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	nios_sys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                                       //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                             //       .reset_req
	);

	nios_sys_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	nios_sys_LCD_ON lcd_on (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (lcd_on_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_on_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_on_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_on_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_on_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_on_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_ON lcd_en (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (lcd_en_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_en_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_en_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_en_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_en_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_en_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_ON lcd_rs (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (lcd_rs_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_rs_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_rs_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_rs_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_rs_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_rs_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_ON lcd_rw (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (lcd_rw_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_rw_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_rw_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_rw_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_rw_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_rw_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA lcd_data (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (lcd_data_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_data_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_data_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_data_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_data_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_data_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led1 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led1_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led2 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led2_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led3 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led3_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led3_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led3_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led3_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led3_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led3_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led4 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led4_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led4_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led4_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led4_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led4_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led4_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led5 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led5_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led5_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led5_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led5_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led5_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led5_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led6 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led6_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led6_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led6_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led6_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led6_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led6_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led7 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led7_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led7_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led7_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led7_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led7_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led7_external_connection_export)                    // external_connection.export
	);

	nios_sys_LCD_DATA led8 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (led8_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led8_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led8_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led8_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led8_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led8_external_connection_export)                    // external_connection.export
	);

	nios_sys_uart_0 uart_0 (
		.clk           (clk_clk),                                                //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address       (uart_0_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_0_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_0_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_0_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_0_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_0_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_0_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                       //                    .dataavailable
		.readyfordata  (),                                                       //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),                         // external_connection.export
		.txd           (uart_0_external_connection_txd),                         //                    .export
		.irq           (irq_mapper_receiver1_irq)                                //                 irq.irq
	);

	nios_sys_switch0 switch0 (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (switch0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch0_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                              //                 irq.irq
	);

	nios_sys_key1 key1 (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address  (key1_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (key1_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (key1_external_connection_export)                  // external_connection.export
	);

	nios_sys_key1 key2 (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address  (key2_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (key2_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (key2_external_connection_export)                  // external_connection.export
	);

	nios_sys_key1 key3 (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address  (key3_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (key3_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (key3_external_connection_export)                  // external_connection.export
	);

	nios_sys_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                              //   irq.irq
	);

	nios_sys_LCD_DATA ledr (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (21),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                      (clk_clk),                                                                            //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_readdatavalid         (),                                                                                   //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (21),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_qsys_0_data_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (17),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led8_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led8_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led8_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led8_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led8_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led8_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led8_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led8_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led8_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led8_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led8_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led8_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led8_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led8_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led8_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led8_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led8_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led7_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led7_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led7_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led7_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led7_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led7_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led7_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led7_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led7_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led7_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led6_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led6_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led6_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led6_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led6_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led6_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led6_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led6_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led6_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led6_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led5_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led4_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led3_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led2_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led1_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (led1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_0_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch0_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (switch0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key3_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (key3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (key3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                   //              (terminated)
		.av_read                  (),                                                                   //              (terminated)
		.av_writedata             (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_chipselect            (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key2_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (key2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (key2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                   //              (terminated)
		.av_read                  (),                                                                   //              (terminated)
		.av_writedata             (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_chipselect            (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key1_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (key1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (key1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                   //              (terminated)
		.av_read                  (),                                                                   //              (terminated)
		.av_writedata             (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_chipselect            (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledr_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_data_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_data_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_data_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_data_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_data_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_data_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_rw_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_rw_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_rw_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_rw_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_rw_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_rw_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_rs_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_rs_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_rs_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_rs_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_rs_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_rs_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_en_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_en_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_en_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_en_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_en_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_en_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_on_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_on_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_on_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_on_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_on_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_on_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_BEGIN_BURST           (76),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.PKT_BURST_TYPE_H          (73),
		.PKT_BURST_TYPE_L          (72),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_THREAD_ID_H           (88),
		.PKT_THREAD_ID_L           (88),
		.PKT_CACHE_H               (95),
		.PKT_CACHE_L               (92),
		.PKT_DATA_SIDEBAND_H       (75),
		.PKT_DATA_SIDEBAND_L       (75),
		.PKT_QOS_H                 (77),
		.PKT_QOS_L                 (77),
		.PKT_ADDR_SIDEBAND_H       (74),
		.PKT_ADDR_SIDEBAND_L       (74),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                     //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                       //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                      //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_BEGIN_BURST           (76),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.PKT_BURST_TYPE_H          (73),
		.PKT_BURST_TYPE_L          (72),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_THREAD_ID_H           (88),
		.PKT_THREAD_ID_L           (88),
		.PKT_CACHE_H               (95),
		.PKT_CACHE_L               (92),
		.PKT_DATA_SIDEBAND_H       (75),
		.PKT_DATA_SIDEBAND_L       (75),
		.PKT_QOS_H                 (77),
		.PKT_QOS_L                 (77),
		.PKT_ADDR_SIDEBAND_H       (74),
		.PKT_ADDR_SIDEBAND_L       (74),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                            //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                           //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                       //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led8_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led8_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led8_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led8_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led8_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led8_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led8_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led8_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led8_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led8_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led8_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led8_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led8_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led8_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led8_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led8_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led8_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                 //                .channel
		.rf_sink_ready           (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led8_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led7_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led7_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led7_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led7_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led7_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led7_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led7_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led7_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                 //                .channel
		.rf_sink_ready           (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led6_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led6_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led6_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led6_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led6_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led6_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led6_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led6_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                 //                .channel
		.rf_sink_ready           (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                 //                .channel
		.rf_sink_ready           (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                 //                .channel
		.rf_sink_ready           (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                 //                .channel
		.rf_sink_ready           (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                 //                .channel
		.rf_sink_ready           (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (led1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                 //                .channel
		.rf_sink_ready           (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_011_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_011_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_011_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_011_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_011_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_011_src_channel),                                                   //                .channel
		.rf_sink_ready           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (switch0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_012_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_012_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_012_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_012_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_012_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_012_src_channel),                                                    //                .channel
		.rf_sink_ready           (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (key3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                 //                .channel
		.rf_sink_ready           (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (key2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_014_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_014_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_014_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_014_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_014_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_014_src_channel),                                                 //                .channel
		.rf_sink_ready           (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (key1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_015_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_015_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_015_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_015_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_015_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_015_src_channel),                                                 //                .channel
		.rf_sink_ready           (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_016_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_016_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_016_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_016_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_016_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_016_src_channel),                                                    //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_017_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_017_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_017_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_017_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_017_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_017_src_channel),                                                 //                .channel
		.rf_sink_ready           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_data_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_data_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                                 //                .channel
		.rf_sink_ready           (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_rw_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                               //                .channel
		.rf_sink_ready           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_rs_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src20_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src20_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src20_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src20_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src20_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src20_channel),                                               //                .channel
		.rf_sink_ready           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_en_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src21_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src21_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src21_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src21_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src21_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src21_channel),                                               //                .channel
		.rf_sink_ready           (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_on_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src22_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src22_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src22_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src22_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src22_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src22_channel),                                               //                .channel
		.rf_sink_ready           (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	nios_sys_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_sys_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	nios_sys_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_sys_id_router id_router_001 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	nios_sys_id_router id_router_002 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                             //          .endofpacket
	);

	nios_sys_id_router id_router_003 (
		.sink_ready         (led8_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led8_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led8_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led8_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led8_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                            //       src.ready
		.src_valid          (id_router_003_src_valid),                                            //          .valid
		.src_data           (id_router_003_src_data),                                             //          .data
		.src_channel        (id_router_003_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_004 (
		.sink_ready         (led7_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led7_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led7_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                            //       src.ready
		.src_valid          (id_router_004_src_valid),                                            //          .valid
		.src_data           (id_router_004_src_data),                                             //          .data
		.src_channel        (id_router_004_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_005 (
		.sink_ready         (led6_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led6_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led6_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                            //       src.ready
		.src_valid          (id_router_005_src_valid),                                            //          .valid
		.src_data           (id_router_005_src_data),                                             //          .data
		.src_channel        (id_router_005_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_006 (
		.sink_ready         (led5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                            //       src.ready
		.src_valid          (id_router_006_src_valid),                                            //          .valid
		.src_data           (id_router_006_src_data),                                             //          .data
		.src_channel        (id_router_006_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_007 (
		.sink_ready         (led4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                            //       src.ready
		.src_valid          (id_router_007_src_valid),                                            //          .valid
		.src_data           (id_router_007_src_data),                                             //          .data
		.src_channel        (id_router_007_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_008 (
		.sink_ready         (led3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                            //       src.ready
		.src_valid          (id_router_008_src_valid),                                            //          .valid
		.src_data           (id_router_008_src_data),                                             //          .data
		.src_channel        (id_router_008_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_009 (
		.sink_ready         (led2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                            //       src.ready
		.src_valid          (id_router_009_src_valid),                                            //          .valid
		.src_data           (id_router_009_src_data),                                             //          .data
		.src_channel        (id_router_009_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_010 (
		.sink_ready         (led1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                            //       src.ready
		.src_valid          (id_router_010_src_valid),                                            //          .valid
		.src_data           (id_router_010_src_data),                                             //          .data
		.src_channel        (id_router_010_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_011 (
		.sink_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                              //       src.ready
		.src_valid          (id_router_011_src_valid),                                              //          .valid
		.src_data           (id_router_011_src_data),                                               //          .data
		.src_channel        (id_router_011_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router id_router_012 (
		.sink_ready         (switch0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                               //       src.ready
		.src_valid          (id_router_012_src_valid),                                               //          .valid
		.src_data           (id_router_012_src_data),                                                //          .data
		.src_channel        (id_router_012_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_id_router id_router_013 (
		.sink_ready         (key3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                            //       src.ready
		.src_valid          (id_router_013_src_valid),                                            //          .valid
		.src_data           (id_router_013_src_data),                                             //          .data
		.src_channel        (id_router_013_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_014 (
		.sink_ready         (key2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                            //       src.ready
		.src_valid          (id_router_014_src_valid),                                            //          .valid
		.src_data           (id_router_014_src_data),                                             //          .data
		.src_channel        (id_router_014_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_015 (
		.sink_ready         (key1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                            //       src.ready
		.src_valid          (id_router_015_src_valid),                                            //          .valid
		.src_data           (id_router_015_src_data),                                             //          .data
		.src_channel        (id_router_015_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_016 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                               //       src.ready
		.src_valid          (id_router_016_src_valid),                                               //          .valid
		.src_data           (id_router_016_src_data),                                                //          .data
		.src_channel        (id_router_016_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_id_router id_router_017 (
		.sink_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                            //       src.ready
		.src_valid          (id_router_017_src_valid),                                            //          .valid
		.src_data           (id_router_017_src_data),                                             //          .data
		.src_channel        (id_router_017_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router_018 id_router_018 (
		.sink_ready         (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                //       src.ready
		.src_valid          (id_router_018_src_valid),                                                //          .valid
		.src_data           (id_router_018_src_data),                                                 //          .data
		.src_channel        (id_router_018_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                           //          .endofpacket
	);

	nios_sys_id_router_018 id_router_019 (
		.sink_ready         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                              //       src.ready
		.src_valid          (id_router_019_src_valid),                                              //          .valid
		.src_data           (id_router_019_src_data),                                               //          .data
		.src_channel        (id_router_019_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router_018 id_router_020 (
		.sink_ready         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                              //       src.ready
		.src_valid          (id_router_020_src_valid),                                              //          .valid
		.src_data           (id_router_020_src_data),                                               //          .data
		.src_channel        (id_router_020_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router_018 id_router_021 (
		.sink_ready         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                              //       src.ready
		.src_valid          (id_router_021_src_valid),                                              //          .valid
		.src_data           (id_router_021_src_data),                                               //          .data
		.src_channel        (id_router_021_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router_018 id_router_022 (
		.sink_ready         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                              //       src.ready
		.src_valid          (id_router_022_src_valid),                                              //          .valid
		.src_data           (id_router_022_src_data),                                               //          .data
		.src_channel        (id_router_022_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                         //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (clk_clk),                            //       clk.clk
		.reset               (rst_controller_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_src_ready),              //      sink.ready
		.sink_channel        (addr_router_src_channel),            //          .channel
		.sink_data           (addr_router_src_data),               //          .data
		.sink_startofpacket  (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_src17_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_006 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src6_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_007 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src7_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src7_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src7_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src7_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src7_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src7_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src7_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src8_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src8_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src8_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src8_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src8_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src8_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src8_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src9_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src9_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src9_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src9_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src9_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src9_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src9_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src9_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_010 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src10_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src10_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src10_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src10_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src10_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src10_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src10_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src10_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_011 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_011_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_011_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_011_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_011_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_011_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_011_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src11_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src11_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src11_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src11_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src11_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src11_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src11_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src11_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_012 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_012_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_012_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_012_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_012_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_012_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_012_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src12_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src12_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src12_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src12_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src12_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src12_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src12_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src12_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_013 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src13_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src13_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src13_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src13_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src13_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src13_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src13_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src13_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_014 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_014_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_014_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_014_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_014_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_014_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_014_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src14_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src14_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src14_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src14_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src14_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src14_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src14_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src14_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_015 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_015_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_015_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_015_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_015_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_015_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_015_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src15_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src15_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src15_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src15_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src15_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src15_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src15_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src15_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_016 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_016_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_016_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_016_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_016_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_016_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_016_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src16_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src16_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src16_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src16_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src16_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src16_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src16_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src16_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_017 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_017_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_017_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_017_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_017_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_017_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_017_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src17_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src17_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src17_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src17_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src17_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src17_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src17_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src17_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_011_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_011_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_012_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_012_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_014_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_014_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_015_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_015_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_016_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_016_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_017_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_017_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_017_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_017_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_017_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_017_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_018 rsp_xbar_demux_018 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_018 rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_018 rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_018 rsp_xbar_demux_021 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_018 rsp_xbar_demux_022 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src1_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src1_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src1_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src1_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src1_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src1_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src1_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src1_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src1_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src1_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src1_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src1_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src1_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src1_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src1_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src1_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src1_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src1_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src1_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src1_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
