library verilog;
use verilog.vl_types.all;
entity lab6_bai1_tb is
end lab6_bai1_tb;
