// nios_sys_tb.v

// Generated using ACDS version 13.0sp1 232 at 2025.04.13.07:59:47

`timescale 1 ps / 1 ps
module nios_sys_tb (
	);

	wire    nios_sys_inst_clk_bfm_clk_clk;       // nios_sys_inst_clk_bfm:clk -> [nios_sys_inst:clk_clk, nios_sys_inst_reset_bfm:clk]
	wire    nios_sys_inst_reset_bfm_reset_reset; // nios_sys_inst_reset_bfm:reset -> nios_sys_inst:reset_reset_n

	nios_sys nios_sys_inst (
		.clk_clk       (nios_sys_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (nios_sys_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_sys_inst_clk_bfm (
		.clk (nios_sys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios_sys_inst_reset_bfm (
		.reset (nios_sys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios_sys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
