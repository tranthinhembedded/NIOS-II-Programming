// nios_sys_tb.v

// Generated using ACDS version 13.0sp1 232 at 2025.04.25.22:56:25

`timescale 1 ps / 1 ps
module nios_sys_tb (
	);

	wire    nios_sys_inst_clk_bfm_clk_clk;       // nios_sys_inst_clk_bfm:clk -> [nios_sys_inst:clk_clk, nios_sys_inst_reset_bfm:clk]
	wire    nios_sys_inst_reset_bfm_reset_reset; // nios_sys_inst_reset_bfm:reset -> nios_sys_inst:reset_reset_n

	nios_sys nios_sys_inst (
		.clk_clk                             (nios_sys_inst_clk_bfm_clk_clk),       //                          clk.clk
		.reset_reset_n                       (nios_sys_inst_reset_bfm_reset_reset), //                        reset.reset_n
		.lcd_data_external_connection_export (),                                    // lcd_data_external_connection.export
		.lcd_rw_external_connection_export   (),                                    //   lcd_rw_external_connection.export
		.lcd_rs_external_connection_export   (),                                    //   lcd_rs_external_connection.export
		.lcd_en_external_connection_export   (),                                    //   lcd_en_external_connection.export
		.lcd_on_external_connection_export   (),                                    //   lcd_on_external_connection.export
		.led8_external_connection_export     (),                                    //     led8_external_connection.export
		.led7_external_connection_export     (),                                    //     led7_external_connection.export
		.led6_external_connection_export     (),                                    //     led6_external_connection.export
		.led5_external_connection_export     (),                                    //     led5_external_connection.export
		.led4_external_connection_export     (),                                    //     led4_external_connection.export
		.led3_external_connection_export     (),                                    //     led3_external_connection.export
		.led2_external_connection_export     (),                                    //     led2_external_connection.export
		.led1_external_connection_export     (),                                    //     led1_external_connection.export
		.uart_0_external_connection_rxd      (),                                    //   uart_0_external_connection.rxd
		.uart_0_external_connection_txd      (),                                    //                             .txd
		.switch0_external_connection_export  (),                                    //  switch0_external_connection.export
		.key3_external_connection_export     (),                                    //     key3_external_connection.export
		.key2_external_connection_export     (),                                    //     key2_external_connection.export
		.key1_external_connection_export     (),                                    //     key1_external_connection.export
		.ledr_external_connection_export     ()                                     //     ledr_external_connection.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_sys_inst_clk_bfm (
		.clk (nios_sys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios_sys_inst_reset_bfm (
		.reset (nios_sys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios_sys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
