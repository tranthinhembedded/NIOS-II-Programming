library verilog;
use verilog.vl_types.all;
entity nios_sys_tb is
end nios_sys_tb;
